module sc_matrix_mult #(

) (
   
);
